//deduplication module
