//selection operator
