//RA controller
