//difference operator
