//Union operator
