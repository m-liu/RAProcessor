//projection operator
