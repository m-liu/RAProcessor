//top BSV file of RA processor
