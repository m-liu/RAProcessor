//cross product operator
