//row marshaller to assemble ddr bursts into table rows
